    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0083;67f8239a;Safari;28E26ABE-48DF-4CE7-B1FB-225F3AAB676A 